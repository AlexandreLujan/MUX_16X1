LIBRARY work;
USE work.MyPackage.all;

ENTITY TestBench IS
END ENTITY;

ARCHITECTURE RTL OF TestBench IS 
	SIGNAL INPUT: BIT_VECTOR(15 DOWNTO 0);
	SIGNAL SE: BIT_VECTOR (3 DOWNTO 0);
	SIGNAL OUTPUT : BIT;
	
BEGIN

	MUX_TEST : MUX_16X1
	port map(
		S => SE(3 downto 0),
		A => INPUT(15 downto 0),
		X => OUTPUT
	);
	
	INPUT <= "1000100010001000" AFTER 0ns, 
				"0100010001000100" AFTER 40ns, 
				"0010001000100010" AFTER 80ns, 
				"0001000100010001" AFTER 120ns; 
   
	SE <= "0000" AFTER 0ns, "1010" AFTER 10ns, "0101" AFTER 20ns, "1111" AFTER 30ns,              
			 "0000" AFTER 40ns, "1010" AFTER 50ns, "0101" AFTER 60ns, "1111" AFTER 70ns,              
			 "0000" AFTER 80ns, "1010" AFTER 90ns, "0101" AFTER 100ns, "1111" AFTER 110ns,              
			 "0000" AFTER 120ns, "1010" AFTER 130ns, "0101" AFTER 140ns, "1111" AFTER 150ns;
	
END ARCHITECTURE;